`ifndef ADDRESSDECODER_V
`define ADDRESSDECODER_V

module AddressDecoder(
    input [15:0] address,
    output reg [2:0] slaveSel
);

    always @(*) begin
        // Default values
        slaveSel = 3'b100;

        // Determine readSelect based on address
        casez (address)
            16'b00??????????????: slaveSel = 3'b001;      // 0x0000 - 0x3FFF
            16'h4000: slaveSel = 3'b010;     // 0x4000
            default: ; // Defaults already set above
        endcase
    end
	 
endmodule
`endif