`timescale 1ns/1ps

module HackComputer_TB;

    // ------------------------------------------------------------------------
    // Parameters
    // ------------------------------------------------------------------------
    localparam integer CLK_PERIOD   = 20;   

    // ------------------------------------------------------------------------
    // UUT interface
    // ------------------------------------------------------------------------
    reg  r_CLK;
    reg  r_RESET_n;

    HackComputer uut (
        .i_CLK      (r_CLK),
        .i_RESET_n  (r_RESET_n)
    );

    // ------------------------------------------------------------------------
    // Clock generation
    // ------------------------------------------------------------------------
    always #(CLK_PERIOD/2) r_CLK = ~r_CLK;

    // ------------------------------------------------------------------------
    // Reset + main stimulus
    // ------------------------------------------------------------------------
    initial begin
        r_CLK       = 1'b0;
        r_RESET_n   = 1'b1;

        // Apply reset
        #(CLK_PERIOD*10);
        r_RESET_n = 1'b0;
        #(CLK_PERIOD*10);
        r_RESET_n = 1'b1;

        // --------------------------------------------------------------------
        repeat (200) @(posedge r_CLK);
        $finish;
    end

    // ------------------------------------------------------------------------
    // VCD dump
    // ------------------------------------------------------------------------
    initial begin
        $display("=== Starting Basic Hack Computer simulation ===");
        $dumpfile("HackComputer_TB.vcd");
        $dumpvars(0, HackComputer_TB);
    end

endmodule
